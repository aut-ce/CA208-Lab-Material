--/*
--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  Designed by Ali Mohammadpour(@alimpk)
--  *******************************************************
--  All Rights reserved (C) 2019-2020
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

-----------------------------------------------------------
---  Module Name: Half Adder
---  Description: Single Bit Half Adder
-----------------------------------------------------------
entity half_adder is
	port (
		a : in  std_logic;
		b : in  std_logic;
		s : out std_logic;
		c : out std_logic
	);
end half_adder;

architecture half_adder_arc of half_adder is
begin

	-- write your code here!

end half_adder_arc;